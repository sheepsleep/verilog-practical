library verilog;
use verilog.vl_types.all;
entity ram_basic_tb is
end ram_basic_tb;
