library verilog;
use verilog.vl_types.all;
entity decode_cmb_tb is
end decode_cmb_tb;
