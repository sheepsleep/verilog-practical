library verilog;
use verilog.vl_types.all;
entity clock_edge_tb is
end clock_edge_tb;
