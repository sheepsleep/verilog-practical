library verilog;
use verilog.vl_types.all;
entity clk_3div_tb is
end clk_3div_tb;
