library verilog;
use verilog.vl_types.all;
entity clk_div_phase_tb is
    generic(
        period          : integer := 5
    );
end clk_div_phase_tb;
